** Library name: gsclib045
** Cell name: DFFSRHQX1
** View name: schematic
.subckt DFFSRHQX1 CK D Q RN SN VDD VSS
*.PININFO  CK:I D:I RN:I SN:I VDD:I VSS:I Q:O
** Above line required by Conformal LEC - DO NOT DELETE

mn26 n20 CKb n21 VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn25 n21 D VSS VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn55 Q qbint VSS VSS g45n1svt L=45e-9 W=260e-9 AD=36.4e-15 AS=36.4e-15 PD=800e-9 PS=800e-9 NRD=538.462e-3 NRS=538.462e-3 M=1
mn35 n30 mout VSS VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn36 n20 CKbb n30 VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn22 RNb RN VSS VSS g45n1svt L=45e-9 W=145e-9 AD=20.3e-15 AS=20.3e-15 PD=570e-9 PS=570e-9 NRD=965.517e-3 NRS=965.517e-3 M=1
mn20 CKb CK VSS VSS g45n1svt L=45e-9 W=145e-9 AD=20.3e-15 AS=20.3e-15 PD=570e-9 PS=570e-9 NRD=965.517e-3 NRS=965.517e-3 M=1
mn45 qbint n35 VSS VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn52 n40 qbint n42 VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn51 n40 RNb n42 VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn32 mout n20 n25 VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn50 n42 SN VSS VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn30 n25 SN VSS VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn40 n35 CKbb mout VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn31 mout RNb n25 VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn21 CKbb CKb VSS VSS g45n1svt L=45e-9 W=145e-9 AD=20.3e-15 AS=20.3e-15 PD=570e-9 PS=570e-9 NRD=965.517e-3 NRS=965.517e-3 M=1
mn53 n35 CKb n40 VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mp26 n20 CKbb n22 VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp25 n22 D VDD VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp52 n43 qbint n41 VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp51 n43 RNb VDD VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp55 Q qbint VDD VDD g45p1svt L=45e-9 W=390e-9 AD=54.6e-15 AS=54.6e-15 PD=1.06e-6 PS=1.06e-6 NRD=358.974e-3 NRS=358.974e-3 M=1
mp36 n20 CKb n31 VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp35 n31 mout VDD VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp32 mout n20 n26 VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp31 n26 RNb VDD VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp22 RNb RN VDD VDD g45p1svt L=45e-9 W=215e-9 AD=30.1e-15 AS=30.1e-15 PD=710e-9 PS=710e-9 NRD=651.163e-3 NRS=651.163e-3 M=1
mp20 CKb CK VDD VDD g45p1svt L=45e-9 W=215e-9 AD=30.1e-15 AS=30.1e-15 PD=710e-9 PS=710e-9 NRD=651.163e-3 NRS=651.163e-3 M=1
mp53 n35 CKbb n41 VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp50 n41 SN VDD VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp45 qbint n35 VDD VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp21 CKbb CKb VDD VDD g45p1svt L=45e-9 W=215e-9 AD=30.1e-15 AS=30.1e-15 PD=710e-9 PS=710e-9 NRD=651.163e-3 NRS=651.163e-3 M=1
mp30 mout SN VDD VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp40 n35 CKb mout VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
.ends DFFSRHQX1
