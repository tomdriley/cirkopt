.MODEL g45n1lvt nmos
.MODEL g45n1svt nmos
.MODEL g45n1hvt nmos
.MODEL g45n2svt nmos
.MODEL g45n1nvt nmos
.MODEL g45n2nvt nmos
.MODEL g45p1lvt pmos
.MODEL g45p1svt pmos
.MODEL g45p1hvt pmos
.MODEL g45p2svt pmos
.MODEL g45p1nvt pmos
.MODEL g45p2nvt pmos


