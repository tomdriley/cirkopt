** Library name: gsclib045
** Cell name: SDFFSRHQX1
** View name: schematic
.subckt SDFFSRHQX1 CK D Q RN SE SI SN VDD VSS
*.PININFO  CK:I D:I RN:I SE:I SI:I SN:I VDD:I VSS:I Q:O
** Above line required by Conformal LEC - DO NOT DELETE

mn13 net534 SI VSS VSS g45n1svt L=45e-9 W=260e-9 AD=36.4e-15 AS=36.4e-15 PD=800e-9 PS=800e-9 NRD=538.462e-3 NRS=538.462e-3 M=1
mn14 Db SE net534 VSS g45n1svt L=45e-9 W=260e-9 AD=36.4e-15 AS=36.4e-15 PD=800e-9 PS=800e-9 NRD=538.462e-3 NRS=538.462e-3 M=1
mn12 Db SEb net522 VSS g45n1svt L=45e-9 W=260e-9 AD=36.4e-15 AS=36.4e-15 PD=800e-9 PS=800e-9 NRD=538.462e-3 NRS=538.462e-3 M=1
mn11 net522 D VSS VSS g45n1svt L=45e-9 W=260e-9 AD=36.4e-15 AS=36.4e-15 PD=800e-9 PS=800e-9 NRD=538.462e-3 NRS=538.462e-3 M=1
mn55 Q qbint VSS VSS g45n1svt L=45e-9 W=260e-9 AD=36.4e-15 AS=36.4e-15 PD=800e-9 PS=800e-9 NRD=538.462e-3 NRS=538.462e-3 M=1
mn35 net514 mout VSS VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn36 n20 CKbb net514 VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn22 RNb RN VSS VSS g45n1svt L=45e-9 W=145e-9 AD=20.3e-15 AS=20.3e-15 PD=570e-9 PS=570e-9 NRD=965.517e-3 NRS=965.517e-3 M=1
mn20 CKb CK VSS VSS g45n1svt L=45e-9 W=145e-9 AD=20.3e-15 AS=20.3e-15 PD=570e-9 PS=570e-9 NRD=965.517e-3 NRS=965.517e-3 M=1
mn45 qbint n35 VSS VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn52 net490 qbint net486 VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn51 net490 RNb net486 VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn50 net486 SN VSS VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn53 n35 CKb net490 VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn10 SEb SE VSS VSS g45n1svt L=45e-9 W=145e-9 AD=20.3e-15 AS=20.3e-15 PD=570e-9 PS=570e-9 NRD=965.517e-3 NRS=965.517e-3 M=1
mn25 Db CKb n20 VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn30 net469 SN VSS VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn32 mout n20 net469 VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn31 mout RNb net469 VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn40 n35 CKbb mout VSS g45n1svt L=45e-9 W=205e-9 AD=28.7e-15 AS=28.7e-15 PD=690e-9 PS=690e-9 NRD=682.927e-3 NRS=682.927e-3 M=1
mn21 CKbb CKb VSS VSS g45n1svt L=45e-9 W=145e-9 AD=20.3e-15 AS=20.3e-15 PD=570e-9 PS=570e-9 NRD=965.517e-3 NRS=965.517e-3 M=1
mp14 Db SEb net453 VDD g45p1svt L=45e-9 W=390e-9 AD=54.6e-15 AS=54.6e-15 PD=1.06e-6 PS=1.06e-6 NRD=358.974e-3 NRS=358.974e-3 M=1
mp13 net453 SI VDD VDD g45p1svt L=45e-9 W=390e-9 AD=54.6e-15 AS=54.6e-15 PD=1.06e-6 PS=1.06e-6 NRD=358.974e-3 NRS=358.974e-3 M=1
mp12 Db SE net445 VDD g45p1svt L=45e-9 W=390e-9 AD=54.6e-15 AS=54.6e-15 PD=1.06e-6 PS=1.06e-6 NRD=358.974e-3 NRS=358.974e-3 M=1
mp11 net445 D VDD VDD g45p1svt L=45e-9 W=390e-9 AD=54.6e-15 AS=54.6e-15 PD=1.06e-6 PS=1.06e-6 NRD=358.974e-3 NRS=358.974e-3 M=1
mp52 net394 qbint net437 VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp51 net437 RNb VDD VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp55 Q qbint VDD VDD g45p1svt L=45e-9 W=390e-9 AD=54.6e-15 AS=54.6e-15 PD=1.06e-6 PS=1.06e-6 NRD=358.974e-3 NRS=358.974e-3 M=1
mp36 n20 CKb net425 VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp35 net425 mout VDD VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp32 mout n20 net417 VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp31 net417 RNb VDD VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp22 RNb RN VDD VDD g45p1svt L=45e-9 W=215e-9 AD=30.1e-15 AS=30.1e-15 PD=710e-9 PS=710e-9 NRD=651.163e-3 NRS=651.163e-3 M=1
mp20 CKb CK VDD VDD g45p1svt L=45e-9 W=215e-9 AD=30.1e-15 AS=30.1e-15 PD=710e-9 PS=710e-9 NRD=651.163e-3 NRS=651.163e-3 M=1
mp53 n35 CKbb net394 VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp50 net394 SN VDD VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp45 qbint n35 VDD VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp25 n20 CKbb Db VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp30 mout SN VDD VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp40 n35 CKb mout VDD g45p1svt L=45e-9 W=310e-9 AD=43.4e-15 AS=43.4e-15 PD=900e-9 PS=900e-9 NRD=451.613e-3 NRS=451.613e-3 M=1
mp21 CKbb CKb VDD VDD g45p1svt L=45e-9 W=215e-9 AD=30.1e-15 AS=30.1e-15 PD=710e-9 PS=710e-9 NRD=651.163e-3 NRS=651.163e-3 M=1
mp10 SEb SE VDD VDD g45p1svt L=45e-9 W=215e-9 AD=30.1e-15 AS=30.1e-15 PD=710e-9 PS=710e-9 NRD=651.163e-3 NRS=651.163e-3 M=1
.ends SDFFSRHQX1
